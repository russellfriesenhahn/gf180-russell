VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vga_clock
  CLASS BLOCK ;
  FOREIGN wrapped_vga_clock ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 288.680 299.000 289.800 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 70.280 299.000 71.400 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.960 296.000 31.080 299.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 164.360 4.000 165.480 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.520 296.000 269.640 299.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 296.000 219.240 299.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 184.520 4.000 185.640 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 50.120 4.000 51.240 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.880 296.000 105.000 299.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.360 1.000 81.480 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 40.040 4.000 41.160 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 268.520 299.000 269.640 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 9.800 299.000 10.920 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.440 296.000 259.560 299.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 208.040 4.000 209.160 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 268.520 4.000 269.640 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 134.120 299.000 135.240 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 29.960 4.000 31.080 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 278.600 4.000 279.720 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.200 296.000 145.320 299.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 278.600 299.000 279.720 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.680 1.000 289.800 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 90.440 299.000 91.560 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.120 296.000 135.240 299.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.520 1.000 185.640 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 154.280 299.000 155.400 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 174.440 4.000 175.560 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.280 1.000 71.400 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 1.000 115.080 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 29.960 299.000 31.080 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.200 4.000 229.320 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.440 296.000 91.560 299.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 103.880 299.000 105.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 164.360 299.000 165.480 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.360 296.000 165.480 299.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 124.040 299.000 125.160 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.440 296.000 175.560 299.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.600 296.000 195.720 299.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.280 296.000 239.400 299.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 298.760 296.000 299.880 299.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 248.360 299.000 249.480 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 1.000 41.160 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.120 296.000 51.240 299.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.120 1.000 135.240 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.440 1.000 175.560 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 258.440 299.000 259.560 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.520 1.000 269.640 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 194.600 299.000 195.720 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.040 296.000 125.160 299.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 144.200 4.000 145.320 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.280 296.000 71.400 299.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.280 296.000 155.400 299.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.280 1.000 239.400 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.440 1.000 91.560 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 80.360 299.000 81.480 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.360 296.000 81.480 299.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 208.040 299.000 209.160 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.880 1.000 21.000 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.600 1.000 279.720 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 60.200 299.000 61.320 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.680 296.000 289.800 299.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.360 4.000 249.480 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.360 1.000 249.480 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.040 1.000 125.160 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 238.280 4.000 239.400 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 228.200 299.000 229.320 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 134.120 4.000 135.240 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 19.880 299.000 21.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 298.760 4.000 299.880 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 296.000 41.160 299.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 194.600 4.000 195.720 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 1.000 219.240 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.960 1.000 31.080 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 124.040 4.000 125.160 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 -0.280 299.000 0.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 174.440 299.000 175.560 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 113.960 299.000 115.080 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.200 1.000 229.320 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 218.120 4.000 219.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 50.120 299.000 51.240 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 154.280 4.000 155.400 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 9.800 4.000 10.920 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 218.120 299.000 219.240 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.440 1.000 259.560 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 238.280 299.000 239.400 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.280 1.000 155.400 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 60.200 4.000 61.320 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 113.960 4.000 115.080 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -0.280 1.000 0.840 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.600 1.000 195.720 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.880 296.000 21.000 299.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 296.000 115.080 299.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.040 296.000 209.160 299.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 19.880 4.000 21.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.120 1.000 51.240 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.800 1.000 10.920 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.360 296.000 249.480 299.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.520 296.000 185.640 299.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.200 1.000 145.320 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.600 296.000 279.720 299.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 40.040 299.000 41.160 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.680 4.000 289.800 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 103.880 4.000 105.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.200 1.000 61.320 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.880 1.000 105.000 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 90.440 4.000 91.560 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 184.520 299.000 185.640 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.360 1.000 165.480 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 70.280 4.000 71.400 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.200 296.000 229.320 299.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.800 296.000 10.920 299.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.200 296.000 61.320 299.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.040 1.000 209.160 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 80.360 4.000 81.480 ;
    END
  END io_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.440 4.000 259.560 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 144.200 299.000 145.320 ;
    END
  END wb_rst_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 282.540 ;
      LAYER Metal2 ;
        RECT 0.700 299.300 298.900 299.510 ;
        RECT 0.700 295.700 9.500 299.300 ;
        RECT 11.220 295.700 19.580 299.300 ;
        RECT 21.300 295.700 29.660 299.300 ;
        RECT 31.380 295.700 39.740 299.300 ;
        RECT 41.460 295.700 49.820 299.300 ;
        RECT 51.540 295.700 59.900 299.300 ;
        RECT 61.620 295.700 69.980 299.300 ;
        RECT 71.700 295.700 80.060 299.300 ;
        RECT 81.780 295.700 90.140 299.300 ;
        RECT 91.860 295.700 103.580 299.300 ;
        RECT 105.300 295.700 113.660 299.300 ;
        RECT 115.380 295.700 123.740 299.300 ;
        RECT 125.460 295.700 133.820 299.300 ;
        RECT 135.540 295.700 143.900 299.300 ;
        RECT 145.620 295.700 153.980 299.300 ;
        RECT 155.700 295.700 164.060 299.300 ;
        RECT 165.780 295.700 174.140 299.300 ;
        RECT 175.860 295.700 184.220 299.300 ;
        RECT 185.940 295.700 194.300 299.300 ;
        RECT 196.020 295.700 207.740 299.300 ;
        RECT 209.460 295.700 217.820 299.300 ;
        RECT 219.540 295.700 227.900 299.300 ;
        RECT 229.620 295.700 237.980 299.300 ;
        RECT 239.700 295.700 248.060 299.300 ;
        RECT 249.780 295.700 258.140 299.300 ;
        RECT 259.860 295.700 268.220 299.300 ;
        RECT 269.940 295.700 278.300 299.300 ;
        RECT 280.020 295.700 288.380 299.300 ;
        RECT 290.100 295.700 298.460 299.300 ;
        RECT 0.700 4.300 298.900 295.700 ;
        RECT 1.140 3.500 9.500 4.300 ;
        RECT 11.220 3.500 19.580 4.300 ;
        RECT 21.300 3.500 29.660 4.300 ;
        RECT 31.380 3.500 39.740 4.300 ;
        RECT 41.460 3.500 49.820 4.300 ;
        RECT 51.540 3.500 59.900 4.300 ;
        RECT 61.620 3.500 69.980 4.300 ;
        RECT 71.700 3.500 80.060 4.300 ;
        RECT 81.780 3.500 90.140 4.300 ;
        RECT 91.860 3.500 103.580 4.300 ;
        RECT 105.300 3.500 113.660 4.300 ;
        RECT 115.380 3.500 123.740 4.300 ;
        RECT 125.460 3.500 133.820 4.300 ;
        RECT 135.540 3.500 143.900 4.300 ;
        RECT 145.620 3.500 153.980 4.300 ;
        RECT 155.700 3.500 164.060 4.300 ;
        RECT 165.780 3.500 174.140 4.300 ;
        RECT 175.860 3.500 184.220 4.300 ;
        RECT 185.940 3.500 194.300 4.300 ;
        RECT 196.020 3.500 207.740 4.300 ;
        RECT 209.460 3.500 217.820 4.300 ;
        RECT 219.540 3.500 227.900 4.300 ;
        RECT 229.620 3.500 237.980 4.300 ;
        RECT 239.700 3.500 248.060 4.300 ;
        RECT 249.780 3.500 258.140 4.300 ;
        RECT 259.860 3.500 268.220 4.300 ;
        RECT 269.940 3.500 278.300 4.300 ;
        RECT 280.020 3.500 288.380 4.300 ;
        RECT 290.100 3.500 298.900 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 298.460 298.950 299.460 ;
        RECT 3.500 290.100 298.950 298.460 ;
        RECT 4.300 288.380 295.700 290.100 ;
        RECT 3.500 280.020 298.950 288.380 ;
        RECT 4.300 278.300 295.700 280.020 ;
        RECT 3.500 269.940 298.950 278.300 ;
        RECT 4.300 268.220 295.700 269.940 ;
        RECT 3.500 259.860 298.950 268.220 ;
        RECT 4.300 258.140 295.700 259.860 ;
        RECT 3.500 249.780 298.950 258.140 ;
        RECT 4.300 248.060 295.700 249.780 ;
        RECT 3.500 239.700 298.950 248.060 ;
        RECT 4.300 237.980 295.700 239.700 ;
        RECT 3.500 229.620 298.950 237.980 ;
        RECT 4.300 227.900 295.700 229.620 ;
        RECT 3.500 219.540 298.950 227.900 ;
        RECT 4.300 217.820 295.700 219.540 ;
        RECT 3.500 209.460 298.950 217.820 ;
        RECT 4.300 207.740 295.700 209.460 ;
        RECT 3.500 196.020 298.950 207.740 ;
        RECT 4.300 194.300 295.700 196.020 ;
        RECT 3.500 185.940 298.950 194.300 ;
        RECT 4.300 184.220 295.700 185.940 ;
        RECT 3.500 175.860 298.950 184.220 ;
        RECT 4.300 174.140 295.700 175.860 ;
        RECT 3.500 165.780 298.950 174.140 ;
        RECT 4.300 164.060 295.700 165.780 ;
        RECT 3.500 155.700 298.950 164.060 ;
        RECT 4.300 153.980 295.700 155.700 ;
        RECT 3.500 145.620 298.950 153.980 ;
        RECT 4.300 143.900 295.700 145.620 ;
        RECT 3.500 135.540 298.950 143.900 ;
        RECT 4.300 133.820 295.700 135.540 ;
        RECT 3.500 125.460 298.950 133.820 ;
        RECT 4.300 123.740 295.700 125.460 ;
        RECT 3.500 115.380 298.950 123.740 ;
        RECT 4.300 113.660 295.700 115.380 ;
        RECT 3.500 105.300 298.950 113.660 ;
        RECT 4.300 103.580 295.700 105.300 ;
        RECT 3.500 91.860 298.950 103.580 ;
        RECT 4.300 90.140 295.700 91.860 ;
        RECT 3.500 81.780 298.950 90.140 ;
        RECT 4.300 80.060 295.700 81.780 ;
        RECT 3.500 71.700 298.950 80.060 ;
        RECT 4.300 69.980 295.700 71.700 ;
        RECT 3.500 61.620 298.950 69.980 ;
        RECT 4.300 59.900 295.700 61.620 ;
        RECT 3.500 51.540 298.950 59.900 ;
        RECT 4.300 49.820 295.700 51.540 ;
        RECT 3.500 41.460 298.950 49.820 ;
        RECT 4.300 39.740 295.700 41.460 ;
        RECT 3.500 31.380 298.950 39.740 ;
        RECT 4.300 29.660 295.700 31.380 ;
        RECT 3.500 21.300 298.950 29.660 ;
        RECT 4.300 19.580 295.700 21.300 ;
        RECT 3.500 11.220 298.950 19.580 ;
        RECT 4.300 9.500 295.700 11.220 ;
        RECT 3.500 1.140 298.950 9.500 ;
        RECT 3.500 0.700 295.700 1.140 ;
      LAYER Metal4 ;
        RECT 59.500 106.490 98.740 217.750 ;
        RECT 100.940 106.490 175.540 217.750 ;
        RECT 177.740 106.490 218.820 217.750 ;
  END
END wrapped_vga_clock
END LIBRARY

