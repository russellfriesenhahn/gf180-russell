VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vga_clock
  CLASS BLOCK ;
  FOREIGN wrapped_vga_clock ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 382.760 399.000 383.880 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 93.800 399.000 94.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 396.000 41.160 399.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 218.120 4.000 219.240 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.880 396.000 357.000 399.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.680 396.000 289.800 399.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 245.000 4.000 246.120 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 66.920 4.000 68.040 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.480 396.000 138.600 399.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.240 1.000 108.360 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 53.480 4.000 54.600 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 355.880 399.000 357.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 13.160 399.000 14.280 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.440 396.000 343.560 399.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 275.240 4.000 276.360 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 355.880 4.000 357.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 177.800 399.000 178.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 40.040 4.000 41.160 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 369.320 4.000 370.440 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.240 396.000 192.360 399.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 369.320 399.000 370.440 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 382.760 1.000 383.880 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 120.680 399.000 121.800 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.800 396.000 178.920 399.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.000 1.000 246.120 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 204.680 399.000 205.800 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 231.560 4.000 232.680 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.800 1.000 94.920 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.920 1.000 152.040 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 40.040 399.000 41.160 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 302.120 4.000 303.240 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.680 396.000 121.800 399.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 137.480 399.000 138.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 218.120 399.000 219.240 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 396.000 219.240 399.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 164.360 399.000 165.480 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.560 396.000 232.680 399.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.440 396.000 259.560 399.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.560 396.000 316.680 399.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.200 396.000 397.320 399.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 329.000 399.000 330.120 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 1.000 54.600 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.920 396.000 68.040 399.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.800 1.000 178.920 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.560 1.000 232.680 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 342.440 399.000 343.560 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.880 1.000 357.000 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 258.440 399.000 259.560 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.360 396.000 165.480 399.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.240 4.000 192.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.800 396.000 94.920 399.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.680 396.000 205.800 399.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.560 1.000 316.680 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.680 1.000 121.800 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 107.240 399.000 108.360 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.240 396.000 108.360 399.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 275.240 399.000 276.360 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.600 1.000 27.720 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.320 1.000 370.440 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 80.360 399.000 81.480 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 382.760 396.000 383.880 399.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 329.000 4.000 330.120 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.000 1.000 330.120 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.360 1.000 165.480 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 315.560 4.000 316.680 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 302.120 399.000 303.240 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 177.800 4.000 178.920 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 26.600 399.000 27.720 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 396.200 4.000 397.320 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 396.000 54.600 399.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.440 4.000 259.560 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.680 1.000 289.800 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 1.000 41.160 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 164.360 4.000 165.480 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 -0.280 399.000 0.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 231.560 399.000 232.680 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 150.920 399.000 152.040 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.120 1.000 303.240 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.680 4.000 289.800 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 66.920 399.000 68.040 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 204.680 4.000 205.800 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 13.160 4.000 14.280 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 288.680 399.000 289.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.440 1.000 343.560 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 315.560 399.000 316.680 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.680 1.000 205.800 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 80.360 4.000 81.480 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 150.920 4.000 152.040 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -0.280 1.000 0.840 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.440 1.000 259.560 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.600 396.000 27.720 399.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.920 396.000 152.040 399.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.240 396.000 276.360 399.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.600 4.000 27.720 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.920 1.000 68.040 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.160 1.000 14.280 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.000 396.000 330.120 399.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.000 396.000 246.120 399.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.240 1.000 192.360 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.320 396.000 370.440 399.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 53.480 399.000 54.600 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 382.760 4.000 383.880 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 137.480 4.000 138.600 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.360 1.000 81.480 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.480 1.000 138.600 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 120.680 4.000 121.800 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 245.000 399.000 246.120 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 1.000 219.240 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 93.800 4.000 94.920 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.120 396.000 303.240 399.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.160 396.000 14.280 399.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.360 396.000 81.480 399.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.240 1.000 276.360 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.240 4.000 108.360 ;
    END
  END io_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 384.460 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 384.460 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 342.440 4.000 343.560 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 191.240 399.000 192.360 ;
    END
  END wb_rst_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 393.120 384.460 ;
      LAYER Metal2 ;
        RECT 0.700 399.300 396.900 399.700 ;
        RECT 0.700 395.700 12.860 399.300 ;
        RECT 14.580 395.700 26.300 399.300 ;
        RECT 28.020 395.700 39.740 399.300 ;
        RECT 41.460 395.700 53.180 399.300 ;
        RECT 54.900 395.700 66.620 399.300 ;
        RECT 68.340 395.700 80.060 399.300 ;
        RECT 81.780 395.700 93.500 399.300 ;
        RECT 95.220 395.700 106.940 399.300 ;
        RECT 108.660 395.700 120.380 399.300 ;
        RECT 122.100 395.700 137.180 399.300 ;
        RECT 138.900 395.700 150.620 399.300 ;
        RECT 152.340 395.700 164.060 399.300 ;
        RECT 165.780 395.700 177.500 399.300 ;
        RECT 179.220 395.700 190.940 399.300 ;
        RECT 192.660 395.700 204.380 399.300 ;
        RECT 206.100 395.700 217.820 399.300 ;
        RECT 219.540 395.700 231.260 399.300 ;
        RECT 232.980 395.700 244.700 399.300 ;
        RECT 246.420 395.700 258.140 399.300 ;
        RECT 259.860 395.700 274.940 399.300 ;
        RECT 276.660 395.700 288.380 399.300 ;
        RECT 290.100 395.700 301.820 399.300 ;
        RECT 303.540 395.700 315.260 399.300 ;
        RECT 316.980 395.700 328.700 399.300 ;
        RECT 330.420 395.700 342.140 399.300 ;
        RECT 343.860 395.700 355.580 399.300 ;
        RECT 357.300 395.700 369.020 399.300 ;
        RECT 370.740 395.700 382.460 399.300 ;
        RECT 384.180 395.700 395.900 399.300 ;
        RECT 0.700 4.300 396.900 395.700 ;
        RECT 1.140 3.500 12.860 4.300 ;
        RECT 14.580 3.500 26.300 4.300 ;
        RECT 28.020 3.500 39.740 4.300 ;
        RECT 41.460 3.500 53.180 4.300 ;
        RECT 54.900 3.500 66.620 4.300 ;
        RECT 68.340 3.500 80.060 4.300 ;
        RECT 81.780 3.500 93.500 4.300 ;
        RECT 95.220 3.500 106.940 4.300 ;
        RECT 108.660 3.500 120.380 4.300 ;
        RECT 122.100 3.500 137.180 4.300 ;
        RECT 138.900 3.500 150.620 4.300 ;
        RECT 152.340 3.500 164.060 4.300 ;
        RECT 165.780 3.500 177.500 4.300 ;
        RECT 179.220 3.500 190.940 4.300 ;
        RECT 192.660 3.500 204.380 4.300 ;
        RECT 206.100 3.500 217.820 4.300 ;
        RECT 219.540 3.500 231.260 4.300 ;
        RECT 232.980 3.500 244.700 4.300 ;
        RECT 246.420 3.500 258.140 4.300 ;
        RECT 259.860 3.500 274.940 4.300 ;
        RECT 276.660 3.500 288.380 4.300 ;
        RECT 290.100 3.500 301.820 4.300 ;
        RECT 303.540 3.500 315.260 4.300 ;
        RECT 316.980 3.500 328.700 4.300 ;
        RECT 330.420 3.500 342.140 4.300 ;
        RECT 343.860 3.500 355.580 4.300 ;
        RECT 357.300 3.500 369.020 4.300 ;
        RECT 370.740 3.500 382.460 4.300 ;
        RECT 384.180 3.500 396.900 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 395.900 399.700 396.340 ;
        RECT 3.500 384.180 399.700 395.900 ;
        RECT 4.300 382.460 395.700 384.180 ;
        RECT 399.300 382.460 399.700 384.180 ;
        RECT 3.500 370.740 399.700 382.460 ;
        RECT 4.300 369.020 395.700 370.740 ;
        RECT 399.300 369.020 399.700 370.740 ;
        RECT 3.500 357.300 399.700 369.020 ;
        RECT 4.300 355.580 395.700 357.300 ;
        RECT 399.300 355.580 399.700 357.300 ;
        RECT 3.500 343.860 399.700 355.580 ;
        RECT 4.300 342.140 395.700 343.860 ;
        RECT 399.300 342.140 399.700 343.860 ;
        RECT 3.500 330.420 399.700 342.140 ;
        RECT 4.300 328.700 395.700 330.420 ;
        RECT 399.300 328.700 399.700 330.420 ;
        RECT 3.500 316.980 399.700 328.700 ;
        RECT 4.300 315.260 395.700 316.980 ;
        RECT 399.300 315.260 399.700 316.980 ;
        RECT 3.500 303.540 399.700 315.260 ;
        RECT 4.300 301.820 395.700 303.540 ;
        RECT 399.300 301.820 399.700 303.540 ;
        RECT 3.500 290.100 399.700 301.820 ;
        RECT 4.300 288.380 395.700 290.100 ;
        RECT 399.300 288.380 399.700 290.100 ;
        RECT 3.500 276.660 399.700 288.380 ;
        RECT 4.300 274.940 395.700 276.660 ;
        RECT 399.300 274.940 399.700 276.660 ;
        RECT 3.500 259.860 399.700 274.940 ;
        RECT 4.300 258.140 395.700 259.860 ;
        RECT 399.300 258.140 399.700 259.860 ;
        RECT 3.500 246.420 399.700 258.140 ;
        RECT 4.300 244.700 395.700 246.420 ;
        RECT 399.300 244.700 399.700 246.420 ;
        RECT 3.500 232.980 399.700 244.700 ;
        RECT 4.300 231.260 395.700 232.980 ;
        RECT 399.300 231.260 399.700 232.980 ;
        RECT 3.500 219.540 399.700 231.260 ;
        RECT 4.300 217.820 395.700 219.540 ;
        RECT 399.300 217.820 399.700 219.540 ;
        RECT 3.500 206.100 399.700 217.820 ;
        RECT 4.300 204.380 395.700 206.100 ;
        RECT 399.300 204.380 399.700 206.100 ;
        RECT 3.500 192.660 399.700 204.380 ;
        RECT 4.300 190.940 395.700 192.660 ;
        RECT 399.300 190.940 399.700 192.660 ;
        RECT 3.500 179.220 399.700 190.940 ;
        RECT 4.300 177.500 395.700 179.220 ;
        RECT 399.300 177.500 399.700 179.220 ;
        RECT 3.500 165.780 399.700 177.500 ;
        RECT 4.300 164.060 395.700 165.780 ;
        RECT 399.300 164.060 399.700 165.780 ;
        RECT 3.500 152.340 399.700 164.060 ;
        RECT 4.300 150.620 395.700 152.340 ;
        RECT 399.300 150.620 399.700 152.340 ;
        RECT 3.500 138.900 399.700 150.620 ;
        RECT 4.300 137.180 395.700 138.900 ;
        RECT 399.300 137.180 399.700 138.900 ;
        RECT 3.500 122.100 399.700 137.180 ;
        RECT 4.300 120.380 395.700 122.100 ;
        RECT 399.300 120.380 399.700 122.100 ;
        RECT 3.500 108.660 399.700 120.380 ;
        RECT 4.300 106.940 395.700 108.660 ;
        RECT 399.300 106.940 399.700 108.660 ;
        RECT 3.500 95.220 399.700 106.940 ;
        RECT 4.300 93.500 395.700 95.220 ;
        RECT 399.300 93.500 399.700 95.220 ;
        RECT 3.500 81.780 399.700 93.500 ;
        RECT 4.300 80.060 395.700 81.780 ;
        RECT 399.300 80.060 399.700 81.780 ;
        RECT 3.500 68.340 399.700 80.060 ;
        RECT 4.300 66.620 395.700 68.340 ;
        RECT 399.300 66.620 399.700 68.340 ;
        RECT 3.500 54.900 399.700 66.620 ;
        RECT 4.300 53.180 395.700 54.900 ;
        RECT 399.300 53.180 399.700 54.900 ;
        RECT 3.500 41.460 399.700 53.180 ;
        RECT 4.300 39.740 395.700 41.460 ;
        RECT 399.300 39.740 399.700 41.460 ;
        RECT 3.500 28.020 399.700 39.740 ;
        RECT 4.300 26.300 395.700 28.020 ;
        RECT 399.300 26.300 399.700 28.020 ;
        RECT 3.500 14.580 399.700 26.300 ;
        RECT 4.300 12.860 395.700 14.580 ;
        RECT 399.300 12.860 399.700 14.580 ;
        RECT 3.500 1.140 399.700 12.860 ;
        RECT 3.500 0.700 395.700 1.140 ;
        RECT 399.300 0.700 399.700 1.140 ;
      LAYER Metal4 ;
        RECT 143.500 60.570 175.540 347.110 ;
        RECT 177.740 60.570 252.340 347.110 ;
        RECT 254.540 60.570 329.140 347.110 ;
        RECT 331.340 60.570 335.860 347.110 ;
  END
END wrapped_vga_clock
END LIBRARY

